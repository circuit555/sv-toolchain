


module foo #(parameter int N = 8) ();
  wire [N-1 : 0] bus;
endmodule;
